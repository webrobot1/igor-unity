<?xml version="1.0" encoding="UTF-8"?><Batch version="2.0"><Options AppVersion="7.5.0"><PathAddFiles><![CDATA[]]></PathAddFiles><PathAddFolder><![CDATA[C:\Users\admin\Desktop\Новая папка (3)\Warrior]]></PathAddFolder></Options><TaskList><Task type="FlipTask" enabled="false"><Horizontal>-1</Horizontal><Vertical>0</Vertical></Task><Task type="CropTask" enabled="true"><Left units="0" base_point="0"><![CDATA[0]]></Left><Right units="0" base_point="2"><![CDATA[0]]></Right><Top units="0" base_point="0"><![CDATA[0]]></Top><Bottom units="0" base_point="2"><![CDATA[0]]></Bottom><Color>#FFFFFF</Color><Alpha>0</Alpha><FillType>0</FillType><Method>1</Method><Width units="1"><![CDATA[66]]></Width><Height units="1"><![CDATA[69]]></Height><Relative>false</Relative><HorizJustification>1</HorizJustification><VertJustification>1</VertJustification></Task><Task type="CropTask" enabled="true"><Left units="0" base_point="0"><![CDATA[0]]></Left><Right units="0" base_point="2"><![CDATA[0]]></Right><Top units="0" base_point="0"><![CDATA[0]]></Top><Bottom units="0" base_point="2"><![CDATA[0]]></Bottom><Color>#FFFFFF</Color><Alpha>0</Alpha><FillType>0</FillType><Method>1</Method><Width units="1"><![CDATA[100]]></Width><Height units="1"><![CDATA[89]]></Height><Relative>false</Relative><HorizJustification>1</HorizJustification><VertJustification>2</VertJustification></Task><Task type="ResizeTask" enabled="true"><Width units="0"><![CDATA[]]></Width><Height units="0"><![CDATA[200]]></Height><DPI><![CDATA[-1]]></DPI><Filter>5</Filter><UseProportions>True</UseProportions><ResizeType>0</ResizeType><ProportionsSize>1</ProportionsSize></Task><Task type="SaveAsTask" enabled="true"><FileName><![CDATA[<Original Name (Without Extension)>]]></FileName><PreserveStruct>True</PreserveStruct><CommonFolder><![CDATA[C:\Users\admin\Desktop\Новая папка (3)\Goblin]]></CommonFolder><FileType></FileType><FilePath><![CDATA[C:\OpenServer\domains\unity\Assets\Resources\Enemy\Goblin\]]></FilePath><FileExists>1</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>95</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed><DDSMIPLevels>8</DDSMIPLevels><DDSMipMapFilter>4</DDSMipMapFilter><DDSFormat>71</DDSFormat><TIFFCompression>0</TIFFCompression><TIFFJPEGColorSpace>2</TIFFJPEGColorSpace><TIFFJPEGQuality>95</TIFFJPEGQuality><TIFFZIPCompression>1</TIFFZIPCompression><TIFFPlanarConf>1</TIFFPlanarConf><DICOMCompression>6</DICOMCompression><DICOMJPEG2000Rate>1</DICOMJPEG2000Rate><DICOMJPEGQuality>95</DICOMJPEGQuality><WEBPLossless>0</WEBPLossless><WEBPQuality>75</WEBPQuality><WEBPMethod>0</WEBPMethod><WEBPTargetSize>0</WEBPTargetSize><WEBPFilterStrength>60</WEBPFilterStrength><WEBPFilterSharpness>0</WEBPFilterSharpness></Task></TaskList></Batch>